module test;

reg[3:0] op;
wire memread;
wire memwrite;
wire branch;
wire alusrc;
wire regdst;
wire regwrite;
wire [1:0] aluop;
wire jump;


endmodule